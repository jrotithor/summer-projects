/*
class class_practice
    int x = 8; 
function return_x()  
	return 8;
endfunction

endclass
*/
module practice(input A, B,C, D, Sel,reset_n, 
input [7:0] v_in,
output [1:0] output2, 
                output [5:0] op_1,
          output out1);
//OSCH #("2.08") osc_int (					
//			.STDBY(1'b0),							
//			.OSC(clk),						
//			.SEDSTDBY());					
		
//string s = "SV";
 logic D1, D2, clk_i;
 clock_counter(.clk_i(clk), .reset_n(reset_n), .clk_o(clk_i));
 mux2(.A(A), .B(B), .Sel(Sel), .Z(D1));
 mux2(.A(C), .B(D), .Sel(Sel), .Z(D2));
 new_adc(.v_in(v_in), .op_1(op_1));
 sv_state_machine(.clk_i(clk_i), .reset_n(reset_n), .in_1(output1), .op_2(output2));
 assign output1 = D1 & D2;
 more_practice(.A(A), .B(B), .out(out1));
endmodule
module mux2(input A, B, Sel,
output reg Z);
 
 always @ *
	 case(Sel)
		 1'b0:	   Z = A;
		 1'b1:     Z = B;
     endcase
endmodule
//typedef struct packed{
//logic [7:0] v_in;


//}v_in;
module new_adc(input [7:0] v_in,
  output [5:0] op_1);
assign op_1 = v_in/4;


endmodule
module sv_state_machine(input clk_i, input [1:0] in_1, input reset_n, 
output logic [1:0] op_2);
parameter S0 = 2'b00;
parameter S1 = 2'b01;
parameter S2 = 2'b10; 
parameter S3 = 2'b11;
logic [1:0]state;
logic [1:0] state_n;
always @ *
	begin
if(in_1 == 2'b00)
	state_n = S1;
else if(in_1 == 2'b01)
	state_n = S2;
else if(in_1 == 2'b10)
	state_n = S3;
else if(in_1 == 2'b11)
	state_n = S0;
else
	state_n = S0;
     end
 always @(posedge clk_i, negedge reset_n)
	begin
if(~reset_n)
	state = S0;
else
	state = state_n;
	     op_2 = state;

end
endmodule

module more_practice(input int A, input int B,
output int out);
struct{

logic [10:0][2:0] a;
logic [10:0][2:0] b;
}types; 
always @ *
	begin
types.a = A;
types.b = B;
  end
int out = A - B;
//$display("%d", out);
 
endmodule    

   module clock_counter(
	input clk_i,		
	input reset_n,
	output logic clk_o
		);
		
		logic [19:0] count;								
														
		
		always @ (posedge clk_i, negedge reset_n)			
			begin
				count <= count + 1;					
				if(!reset_n)
					begin
						clk_o <= 0;
						count <= 0;						
					end
				else
					if(count >=86666)					
						begin							
							clk_o <= ~clk_o;	
							count <= 0;					
						end
			end 
		  
		
endmodule

// TOOL:     vlog2tf
// DATE:     Mon May 11 18:48:09 2015
 
// TITLE:    Lattice Semiconductor Corporation
// MODULE:   Clock_source
// DESIGN:   Clock_source
// FILENAME: Clock_source_tf.v
// PROJECT:  Unknown
// VERSION:  2.0
// This file is auto generated by the Diamond


`timescale 1 ms / 1 ms

// Define Module for Test Fixture

// TOOL:     vlog2tf
// DATE:     Mon May 11 18:48:09 2015
 
// TITLE:    Lattice Semiconductor Corporation
// MODULE:   Clock_source
// DESIGN:   Clock_source
// FILENAME: Clock_source_tf.v
// PROJECT:  Unknown
// VERSION:  2.0
// This file is auto generated by the Diamond


`timescale 1 ms / 1 ms

// Define Module for Test Fixture
module practice_tf();
 
// Inputs
    logic A;
	logic B;
	logic C;
	logic D;
	logic Sel;
	logic reset_n;
	logic [7:0] v_in;
	


// Outputs
 logic [1:0]output2;   
  logic [5:0] op_1;
    logic out1;
   


// Bidirs


// Instantiate the UUT
// Please check and add your parameters manually
    practice UUT (
        .A(A), 
        .B(B), 
        .C(C), 
        .D(D), 
        .Sel(Sel), 
        .reset_n(reset_n), 
        .v_in(v_in),
		.output2(output2),
		.op_1(op_1),
		.out1(out1)
        );


// Initialize Inputs
// You can add your stimulus here
    initial begin
       $dumpfile("dump.vcd");
  $dumpvars(1,practice_tf);
          reset_n = 0; A = 0; B = 0; C = 0; D = 0; Sel = 0; v_in = 0;
		  #10 reset_n = 1; A = 1; B = 1;
      	  #10 v_in = 125;
          #10 C = 1;
      	  #10 D = 1;
	
	
	
    end

endmodule // Clock_source_tf
